library ieee;
use ieee.std_logic_1164.ALL;
use ieee.std_logic_unsigned.ALL;
use ieee.numeric_std.ALL;

entity down_dec is
	port (Data_in : in std_logic_vector(23 downto 0);
			Data_out_I : out std_logic_vector(23 downto 0);
			Data_out_Q : out std_logic_vector(23 downto 0);
			clk_in : in std_logic; 
			clk_sample : in std_logic; 
			rx_att : in std_logic_vector(1 downto 0);
			clk_out : out std_logic
			);
end down_dec;

architecture down_dec_arch of down_dec is
	
type longbuffer is array (649 downto 0) of signed (23 downto 0);
type filt_type is array (319 downto 0) of signed (23 downto 0);

signal Ia : longbuffer;
signal Qa : longbuffer;
	 
constant filtkoeff : filt_type :=

-- Scilab:
-->[v,a,f] = wfir ('lp', 640, [25/625 0], 'hn', 0);
-->round(v*2^ 26)

	("000000000000000000000000",
    "111111111111111111111110",
    "111111111111111111111010",
    "111111111111111111110100",
    "111111111111111111101110",
    "111111111111111111101100",
    "111111111111111111110001",
    "000000000000000000000000",
    "000000000000000000011010",
    "000000000000000001000001",
    "000000000000000001110010",
    "000000000000000010101011",
    "000000000000000011100110",
    "000000000000000100011100",
    "000000000000000101000101",
    "000000000000000101011001",
    "000000000000000101001111",
    "000000000000000100100001",
    "000000000000000011001100",
    "000000000000000001001110",
    "111111111111111110101010",
    "111111111111111011101000",
    "111111111111111000010100",
    "111111111111110100111101",
    "111111111111110001110110",
    "111111111111101111010001",
    "111111111111101101100100",
    "111111111111101100111111",
    "111111111111101101110011",
    "111111111111110000001000",
    "111111111111110100000000",
    "111111111111111001011000",
    "000000000000000000000000",
    "000000000000000111100100",
    "000000000000001111100110",
    "000000000000010111100011",
    "000000000000011110110100",
    "000000000000100100110010",
    "000000000000101000110101",
    "000000000000101010011101",
    "000000000000101001010000",
    "000000000000100101000001",
    "000000000000011101101110",
    "000000000000010011100100",
    "000000000000000111000000",
    "111111111111111000101010",
    "111111111111101001011010",
    "111111111111011010001111",
    "111111111111001100001110",
    "111111111111000000011101",
    "111111111110110111111101",
    "111111111110110011101000",
    "111111111110110100000111",
    "111111111110111001110100",
    "111111111111000100110000",
    "111111111111010100101000",
    "111111111111101000101110",
    "000000000000000000000000",
    "000000000000011001001000",
    "000000000000110010100000",
    "000000000001001010011011",
    "000000000001011111001001",
    "000000000001101111000010",
    "000000000001111000101010",
    "000000000001111010111010",
    "000000000001110101000111",
    "000000000001100111001000",
    "000000000001010001010011",
    "000000000000110100100110",
    "000000000000010010011111",
    "111111111111101100111010",
    "111111111111000110001010",
    "111111111110100000110000",
    "111111111101111111010010",
    "111111111101100100001111",
    "111111111101010001110011",
    "111111111101001001101111",
    "111111111101001101001101",
    "111111111101011100101001",
    "111111111101110111110000",
    "111111111110011101011001",
    "111111111111001011101010",
    "000000000000000000000000",
    "000000000000110111010001",
    "000000000001101101111111",
    "000000000010100000011111",
    "000000000011001011001101",
    "000000000011101010111011",
    "000000000011111100111101",
    "000000000011111111011001",
    "000000000011110001010001",
    "000000000011010010101001",
    "000000000010100100101110",
    "000000000001101001101110",
    "000000000000100100111000",
    "111111111111011010001110",
    "111111111110001110010111",
    "111111111101000110001110",
    "111111111100000110101100",
    "111111111011010100010111",
    "111111111010110011001000",
    "111111111010100101111111",
    "111111111010101110101111",
    "111111111011001101110010",
    "111111111100000010001001",
    "111111111101001001010111",
    "111111111110011111101000",
    "000000000000000000000000",
    "000000000001100100101000",
    "000000000011000111001010",
    "000000000100100001000100",
    "000000000101101100001000",
    "000000000110100010110100",
    "000000000111000000101110",
    "000000000111000010110110",
    "000000000110100111111000",
    "000000000101110000010111",
    "000000000100011110101111",
    "000000000010110111001101",
    "000000000000111111101000",
    "111111111110111111000110",
    "111111111100111101100110",
    "111111111011000011011111",
    "111111111001011000111110",
    "111111111000000101100100",
    "111111110111001111100110",
    "111111110110111011101011",
    "111111110111001100011100",
    "111111111000000010001100",
    "111111111001011010111000",
    "111111111011010010000101",
    "111111111101100001001111",
    "000000000000000000000000",
    "000000000010100100101011",
    "000000000101000100110110",
    "000000000111010101111111",
    "000000001001001110001100",
    "000000001010100100110001",
    "000000001011010010111010",
    "000000001011010100001100",
    "000000001010100110111010",
    "000000001001001100010100",
    "000000000111001000101011",
    "000000000100100011000000",
    "000000000001100100110011",
    "111111111110011001011101",
    "111111111011001101101001",
    "111111111000001110011101",
    "111111110101101000101010",
    "111111110011100111110011",
    "111111110010010101011100",
    "111111110001111000011110",
    "111111110010010100100100",
    "111111110011101001110110",
    "111111110101110100101111",
    "111111111000101110000101",
    "111111111100001011100001",
    "000000000000000000000000",
    "000000000011111100100100",
    "000000000111110001001111",
    "000000001011001110000000",
    "000000001110000011111011",
    "000000010000000110000010",
    "000000010001001010010001",
    "000000010001001010010000",
    "000000010000000011110011",
    "000000001101111001001010",
    "000000001010110001000011",
    "000000000110110110011000",
    "000000000010010111100111",
    "111111111101100110000001",
    "111111111000110100101000",
    "111111110100010111000011",
    "111111110000100000001111",
    "111111101101100001001111",
    "111111101011101000000100",
    "111111101010111110101010",
    "111111101011101010001011",
    "111111101101101010011101",
    "111111110000111001111010",
    "111111110101001101101011",
    "111111111010010110001100",
    "000000000000000000000000",
    "000000000101110100111101",
    "000000001011011101011111",
    "000000010000100010000110",
    "000000010100101100111001",
    "000000010111101011000001",
    "000000011001001101111011",
    "000000011001001100100000",
    "000000010111100011110010",
    "000000010100010111010111",
    "000000001111110001010001",
    "000000001010000001100111",
    "000000000011011101101111",
    "111111111100011110111011",
    "111111110101100000111110",
    "111111101111000000011101",
    "111111101001011000111100",
    "111111100101000011001001",
    "111111100010010011010110",
    "111111100001010111110111",
    "111111100010011000000011",
    "111111100101010011100000",
    "111111101010000001111111",
    "111111110000010011101000",
    "111111110111110001101110",
    "000000000000000000000000",
    "000000001000011110010001",
    "000000010000101010010100",
    "000000011000000010000101",
    "000000011110000101110010",
    "000000100010011010000100",
    "000000100100101001111000",
    "000000100100100111111101",
    "000000100010001111111110",
    "000000011101100111000100",
    "000000010110111011101111",
    "000000001110100101010011",
    "000000000101000010101000",
    "111111111010111000011010",
    "111111110000101110111110",
    "111111100111001111110110",
    "111111011111000011001010",
    "111111011000101101000001",
    "111111010100101011000111",
    "111111010011010010100101",
    "111111010100101110011001",
    "111111011000111110011011",
    "111111011111110111000001",
    "111111101001000001011000",
    "111111110011111100101110",
    "000000000000000000000000",
    "000000001100011100010001",
    "000000011000011111011110",
    "000000100011010111100000",
    "000000101100010101011110",
    "000000110010110000101011",
    "000000110110001001011100",
    "000000110110001011011110",
    "000000110010101111011100",
    "000000101011111011111010",
    "000000100010000101011000",
    "000000010101101101011101",
    "000000000111100001001011",
    "111111111000010110100001",
    "111111101001001001010000",
    "111111011010110111011110",
    "111111001110011101100110",
    "111111000100110010100101",
    "111110111110100100010000",
    "111110111100010100000010",
    "111110111110010100011011",
    "111111000100100111010010",
    "111111001110111101001000",
    "111111011100110101011100",
    "111111101101100000001001",
    "000000000000000000000000",
    "000000010011001110000001",
    "000000100101111101100000",
    "000000110111000000101110",
    "000001000101001101101101",
    "000001001111100011000100",
    "000001010101001100011110",
    "000001010101100110011000",
    "000001010000100000111111",
    "000001000110000010000100",
    "000000110110100101011010",
    "000000100010111100000111",
    "000000001100001010010110",
    "111111110011100011111110",
    "111111011010100111111100",
    "111111000010111010111100",
    "111110101110000001011001",
    "111110011101011001001001",
    "111110010010010011011011",
    "111110001101101111001010",
    "111110010000010100010011",
    "111110011010010000000111",
    "111110101011010011001100",
    "111111000010110000110100",
    "111111011111100000010101",
    "000000000000000000000000",
    "000000100010011001101100",
    "000001000100101000111001",
    "000001100100100001111110",
    "000001111111111010001100",
    "000010010100110000000001",
    "000010100001010011011011",
    "000010100100001101100111",
    "000010011100100111101010",
    "000010001010001111101101",
    "000001101101011100011100",
    "000001000111001110010101",
    "000000011001001110110110",
    "111111100101101101001100",
    "111110101111011000111111",
    "111101111001011010111000",
    "111101000111001011011111",
    "111100011100001001001001",
    "111011111011101100101110",
    "111011101000111110011010",
    "111011100110101010101111",
    "111011110110111000100100",
    "111100011011000000100111",
    "111101010011100110111001",
    "111110100000010110011110",
    "000000000000000000000000",
    "000001110000011010110110",
    "000011101110101001001000",
    "000101110110111110011001",
    "001000000101001000101000",
    "001010010100011011010011",
    "001100011111111011111010",
    "001110100010101111010110",
    "010000011000000111100111",
    "010001111011110001000011",
    "010011001001111110101011",
    "010011111111110100101100",
    "010100011011010000111110"
	);

--attribute ramstyle : string;
--attribute ramstyle of filtkoeff : constant is "M4K";

signal sample : boolean := false;
signal sampled : boolean := false;

signal I_asynch,Q_asynch, I_synch, Q_synch : signed (23 downto 0);

signal filtk : signed(23 downto 0);
signal prod_I : signed (47 downto 0);
signal prod_Q : signed (47 downto 0);
signal mac_I : signed (65 downto 0);
signal mac_Q : signed (65 downto 0);

signal write_pointer, write_pointer_last : integer range 0 to 649 := 600;
signal read_pointer : integer range 0 to 649;
signal clk_out_next : boolean := false;

signal inbuffer : signed(23 downto 0);
	
begin

downconversion : process (clk_in)
	variable ns : integer range 0 to 3 := 0;	
	begin	
		if clk_in'event and clk_in = '1' then		
			if clk_out_next = true then
				clk_out <= '1';
			else
				clk_out <= '0';
			end if;

			if sample = true then
				sampled <= true;			
			elsif sampled = true then
				if ns = 0 then
					Ia(write_pointer) <= inbuffer;  				-- 1
					Qa(write_pointer) <= to_signed(0,24); 		-- 0
					ns := 1;
				elsif ns = 1 then
					Ia(write_pointer) <= to_signed(0,24);		-- 0
					Qa(write_pointer) <= inbuffer;			-- 1
					ns := 2;
				elsif ns = 2 then
					Ia(write_pointer) <= (not inbuffer) + 1; -- -1
					Qa(write_pointer) <= to_signed(0,24); 	 -- 0
					ns := 3;
				elsif ns = 3 then
					Ia(write_pointer) <= to_signed(0,24);		-- 0
					Qa(write_pointer) <= (not inbuffer) + 1; -- -1
					ns := 0;
				end if;		
				write_pointer_last <= write_pointer;
				sampled <= false;
				if write_pointer = 0 or write_pointer > 649 then
					write_pointer <= 649;
				else
					write_pointer <= write_pointer - 1;
				end if;	
			end if;
			I_asynch <= Ia(read_pointer);
			Q_asynch <= Qa(read_pointer);
			I_synch <= I_asynch;
			Q_synch <= Q_asynch;
		end if;
	end process;
	
filter : process (clk_in)
	variable n : integer range 0 to 649 := 0;
	variable nn : integer range 0 to 319;
	variable m : integer range 0 to 8 := 0;
	variable filter_start_pointer : integer range 0 to 649 := 100;
	variable p : integer range 0 to 1500;

	begin	
		if clk_in'event and clk_in = '1' then
			if sampled = true then		
				if m = 7 then  -- start filtering every 8 samples
					clk_out_next <= true;
					filter_start_pointer := write_pointer_last;
					m := 0;    -- written samples
					n := 0;	  -- multiplication steps						
					prod_I <= to_signed(0,48);
					prod_Q <= to_signed(0,48);	
					mac_I <= to_signed(0,66);
					mac_Q <= to_signed(0,66);	
					filtk <= filtkoeff(0);
				else
					clk_out_next <= false;
					m := m + 1;
				end if;
			end if;
			
			p := filter_start_pointer + n;
			if p > 649 then
				read_pointer <= p - 650;
			else
				read_pointer <= p;
			end if;
					
			if n > 2 and n < 642 then  -- valid data after two reads
				if n < 322 then
					nn := n - 2;   -- nn = 1 to 319
				else 
					nn := 641 - n; -- nn = 319 to 0, symmetric filter, only half of the taps need to be stored
				end if;
				filtk <= filtkoeff(nn);
            prod_I <= I_synch*filtk; 
				prod_Q <= Q_synch*filtk;
				mac_I <= mac_I + prod_I;
				mac_Q <= mac_Q + prod_Q;
				n := n + 1;
			elsif n = 642 then
				prod_I <= I_synch*filtk; 
				prod_Q <= Q_synch*filtk;
				mac_I <= mac_I + prod_I;
				mac_Q <= mac_Q + prod_Q;
				n := n + 1;
			elsif n = 643 then
				mac_I <= mac_I + prod_I;
				mac_Q <= mac_Q + prod_Q;
				n := n + 1;
			elsif n = 644 then
				if rx_att = "11" then
					Data_out_I <= std_logic_vector(mac_I + to_signed(67108864,66))(50 downto 27);  
					Data_out_Q <= std_logic_vector(mac_Q + to_signed(67108864,66))(50 downto 27);
				elsif rx_att = "10" then
					Data_out_I <= std_logic_vector(mac_I + to_signed(33554432,66))(49 downto 26); 
					Data_out_Q <= std_logic_vector(mac_Q + to_signed(33554432,66))(49 downto 26);
				elsif rx_att = "01" then
					Data_out_I <= std_logic_vector(mac_I + to_signed(16777216,66))(48 downto 25);  
					Data_out_Q <= std_logic_vector(mac_Q + to_signed(16777216,66))(48 downto 25);
				else
					Data_out_I <= std_logic_vector(mac_I + to_signed(8388608,66))(47 downto 24);  
					Data_out_Q <= std_logic_vector(mac_Q + to_signed(8388608,66))(47 downto 24);
				end if;				
			else
            n := n + 1;
         end if;
			
		end if;
	end process;
	
	
	sample_ff : process(clk_sample, sampled)
	begin
		if sampled = true then
			sample <= false;
		elsif clk_sample'event and clk_sample = '1' then
			inbuffer <= signed(data_in);
			sample <= true;
		end if;
	end process;
	
	
end down_dec_arch;