library ieee;
use ieee.std_logic_1164.ALL;
--use ieee.std_logic_unsigned.ALL;
use ieee.numeric_std.ALL;

entity audio_synch is
	port (
			audio_in : in std_logic_vector(15 downto 0);
			codec_clk : in std_logic;
			i2s_clk : in std_logic;
			audio_out : out std_logic_vector(15 downto 0)
			);
end audio_synch;

architecture arch of audio_synch is

signal in_reg_1 : std_logic_vector(15 downto 0);

begin

sample : process(codec_clk)
	begin
		if codec_clk'event and codec_clk = '1' then
			in_reg_1 <= audio_in;
		end if;
	end process;

sample_i2s : process(i2s_clk)
	begin
		if i2s_clk'event and i2s_clk = '1' then
			audio_out <= in_reg_1;
		end if;
	end process;

end arch;




library ieee;
use ieee.std_logic_1164.ALL;
--use ieee.std_logic_unsigned.ALL;
use ieee.numeric_std.ALL;

entity i2s_master is
	port (clk0 : in std_logic;
			sample_clk : in std_logic;
			I_data_in : in std_logic_vector(23 downto 0);
			Q_data_in : in std_logic_vector(23 downto 0);
			iqswap : in std_logic;
			audio_out_l : out std_logic_vector(15 downto 0);
			audio_out_r : out std_logic_vector(15 downto 0);
			audio_in : in std_logic_vector(15 downto 0);
			bclk : buffer std_logic;
			lrclk : out std_logic;
			dout : out std_logic;
			din : in std_logic;
			tx : in std_logic;
			key : in std_logic;
			loopback : in std_logic
			);
end i2s_master;

architecture arch of i2s_master is

signal data_reg_1, data_reg_2 : std_logic_vector(31 downto 0);
signal receive_reg, data_received_r, data_received_l : std_logic_vector(31 downto 0);
signal sample : std_logic;
signal sample_rst : std_logic;
signal clockdiv : integer range 0 to 21;
 
begin

	dout <= data_reg_2(31);   --  ändra till process för att ge 96 kHz
	--bclk <= clockdiv(1);
	
	audio_out_l <= data_received_l (31 downto 16);
	audio_out_r <= data_received_r (31 downto 16);
	
	clockdivider : process(clk0)
	begin
		if clk0'event and clk0 = '1' then
			if clockdiv = 20 then
				bclk <= not bclk;
				clockdiv <= 0;
			else
				clockdiv <= clockdiv + 1;
			end if;
		end if;
	end process;
		
	sample_ff : process(sample_rst,sample_clk)
	begin
		if sample_rst = '1' then
			sample <= '0';
		elsif sample_clk'event and sample_clk = '1' then
			sample <= '1';
		end if;
	end process;

	bitclk : process(bclk)
	variable bitcount : integer range 0 to 63;
	begin
		if bclk'event and bclk = '0' then
			if sample = '1' then
				if tx = '1' then
					if loopback = '0' then
						data_reg_1 <= audio_in & "000000000000000" & key;
					else
						data_reg_1 <= data_received_l(31 downto 1) & key;
					end if;
				elsif iqswap = '0' then
					data_reg_1 <= I_data_in & "00000000";
				else
					data_reg_1 <= Q_data_in & "00000000";
				end if;
				sample_rst <= '1';
				bitcount := 63;
				lrclk <= '0';
				data_reg_2 <= data_reg_2(30 downto 0) & '0';
			elsif bitcount = 63 then
				bitcount := 0;
				data_reg_2 <= data_reg_1;
				sample_rst <= '0';
				data_received_r <= receive_reg;
			elsif bitcount = 30 then
				lrclk <= '1';
				bitcount := 31;
				if tx = '1' then
					if loopback = '0' then
						data_reg_1 <= audio_in & "000000000000000" & key;
					else
						data_reg_1 <= data_received_r(31 downto 1) & key;
					end if;
				elsif iqswap = '0' then
					data_reg_1 <= Q_data_in & "00000000";
				else
					data_reg_1 <= I_data_in & "00000000";
				end if;
				data_reg_2 <= data_reg_2(30 downto 0) & '0';
			elsif bitcount = 31 then
				bitcount := 32;
				data_reg_2 <= data_reg_1;
				data_received_l <= receive_reg;
			else
				bitcount := bitcount + 1;
				data_reg_2 <= data_reg_2(30 downto 0) & '0';
			end if;
		elsif bclk'event and bclk = '1' then
			receive_reg <= receive_reg(30 downto 0) & din;
		end if;
	end process;

end arch;